`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.07.2025 13:02:46
// Design Name: 
// Module Name: class_top_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module class_top_tb;
    reg clk;
    reg [1:0]prst;
    reg [19:0]model_params;
    reg [14:0]count = 0;
    reg [511:0] total_img;
    reg tvalid;
    reg [7:0]bram_addr_a;
    reg [3:0]bram_addr_a2;
    reg [3:0]label;
    reg [3:0]calc_label;
    reg [181:0]clause_write;
    reg [1259:0]weight_write;
    reg [10:0] success;
    reg [10:0] fail;
    reg opm;
    wire [4:0]output_params;
    wire tready;
    
     initial clk = 1;
    always #5 clk = ~clk;
    integer img_count = 0;
    class_top
    uut
    (clk,prst,model_params,total_img,tvalid,img_count,bram_addr_a,bram_addr_a2,clause_write,weight_write,tready,output_params);
    initial 
    begin    
        count = 0;
        success = 0;
        fail = 0; 
        prst = 3;
        model_params = 20'b1010_010001100_001_1_111;
        #20
        prst = 0;
        tvalid = 1;
        #10
//number 0
       total_img = 512'b00000000000000011100000001100000000000000001100000000110000000000000000110000000011000000000000000011000000001100000000000000001100000000110000000000000000110000000111000000000000000011000000011100000000000000001110000001110000000000000000111000001110000000000000000001100000111000000000000000000111100011100000000000000000001111111110000000000000000000111111110000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10
       total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000011111111000000000000000000011111011110000000000000000001110000111000000000000000001110000001100000000000000000110000000110;
       
        #10        
        bram_addr_a2 = 0;
        weight_write = 0;
        #10 
        weight_write = 1260'b001011101000000000100000000011000100110100000100101100000000000000000000000011010000111110111111110111110010010101110111111101010000101000000000100000000001110100000010000100000000000000000010001111000000010000000000000000000111000000010011000000000000000000000111101100010001000000000000000000000110010011100000000000000000100000000000000000000000000000000000000011011010001110000000000100000000110011010000000000011010110100000000000000000000000000000000000001011110001101100000000000000110101000000000100011101000000100011000110000000000100000000011111011100000000010010110110110001000110010000000000000100001100000000011111111111111100000000000000111110100000000000000000000010011110001111110101011000000000010010111000011011011001100000000000010000000000101101001011010000000000111111010000000000000000100000000000100000000000000000011010001000000000110100110011001101011100000010110001001100100000000000011000110000000000000101000001111001011011010000000000111101110011100010100000000000110101100000000000000000000000000010100010100000000111111011001101000101100111010011101000000000000110001000000000111101111011100100010110110100000000000000000110110010010111110101000001000010100010001001000000000000000000000000000000000000111110000100000000100000000; 
        #10 
        bram_addr_a2 = 1;
        weight_write = 1260'b001010000110101011110100110100000000111011111000000000000000000100000000000000000000100101000000100100000000000101100000000011000000000000000000000000000010010010110011101100000000000000000100000000001011101000000000000000000001101110000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000100000000100000000000000000000000000111011000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010001110110011100000000000101001111000000000010111011000000110000000000000000000000000000000000000100000000101011111100000000111110111000000000000100011001010010000000000000001111000000000001010100100000000000000000000000000010100100000000000000000000000000000111110100000000000000000000001000000100000000100000000000000000100000000000000000111111010000000000000000000000000000000000000001000111001100011001100000000000000000000000100000000000000000000000000000000000010001001100000000000000000000000000000000000100000000100000000011001110000000000111001011000000000100000000011000011000000001100000000010101000100000000000000000111101101000000000000001011000000000000000000000000000011010000000000000000000000000000000111010010000000000000000000000000000100000000000000000000000000000000000111110001; 
        #10 
        bram_addr_a2 = 2;
        weight_write = 1260'b001000001011011000100000000100000000111011111100000000000000000000000000001000010001000101000000100110110110010011011000000000001010111000000000000111010001001101001000101100000000001010101111010001111100101011110001000000000111011110111011001000000000000000000001100001100000000000000000000000000000010110001100001011111111001010100001001010011111010000000000000011011000000000000000000010100000010011000001110001100000000010110011000000000000101101000000000010001110001101110000000000000011101000000000111011101000000110000000000000000000011000101000000000010000001111001110010000000101001000000000000111101010111111001000000000100000000000000000110111101010001111011010011000000000100000000010111111000000000001011001111101000000001100000000000100000000111100101111111110011111100001001100000000000000000110000000000100000000000000000111111110101110010000101010000000000111110010000000000101111100000000000111000111011110011111010111110111000100000000000000000101001000100000000001000001110110100011100111100000000000000000000011111000101001000000001110011011100010000001000100000000000000110100000000000111111001000000000010011111010010011100000000111001110011011101000111100000001111001011000000000000000000000100000000000000000111001011011101011100000000; 
         #10 
        bram_addr_a2 = 3;
        weight_write = 1260'b101100000000100110110100110100000000010111100001111010000000000010001011001111011111110010000000100010001110111110111111110110010010101000000000100000000010001110001001101101000110010111000110111000111011001011000110000000000100000000010011101000000000000000000001010011100000000000000000000000000010001011010100101000000000100000000000010101100000000011111111000011110010001110000000000101010001000010000000000000100000000100000000000000000011101010011111111000000000001101010000000000000011001000000000100000000111111110000000000011000110100000000000000000001001110101011111100000000101001000000000000101000100111000101000000000000011110000000000100000000100000000010110101000000000000000000010111111011100011100110101111101100010011110000000000100000000010101011010011111000000000001000000000000000000000100000000000111110110011110001000110000000000000000000101000000000010000111000000000010010101000000000000000000100000000000000000000111010100110011000000000110000101100000000001001000000000000100000000100000001000000000010010001101000101000000001100000000100000000001101101000000000000101100000000000111111111000000000110110100111111101000000000100000000101001000101110101111100110100000000011110001000000000100001010000000000011000010000000000000000000; 
         #10 
        bram_addr_a2 = 4;
        weight_write = 1260'b111111011001100011000111011001101101000101110001111101000000000001010111100000000111111010111110100100000000001000000000000011100000000011111111010110101100000000100000100001100001001010101100011010111010011000000000000000000000111001100000000000000000000000000001001011010001000011111111000000000100000000000010111000000000100000000010000110000000000000000000111001111001011110000000000100000000100000000011000110001111110000000000011111111100000000000000000000000000100000000000000000101111100000000000100000000000000100000000000000000000000000000000000000100000000000000000100000000101001000011111111000100001110011001000000000000010101011111000100110111100000000100000000001111101000101101000000000000000000111110111000011110000000000000000000000101110100000000001010100000000000000110011000000000111100011000000000001010101000000000000000000001000111111100000010011100010000111011010101100000000000000000100011101000000000011101011110111000100000000000000000000000000101110101001111010100000000000111011011001010000000000100000000000101001000000001000100111010001101100000000000000000111110101000000000000001011010110011100000000010011111001001010000000000000000000101110101111101010010100110000000000000000000001111101000000000100000000100000000010010111; 
         #10 
        bram_addr_a2 = 5;
        weight_write = 1260'b100000000000000000110100110110011110100000000000011100000000000010101001000001101111110110000000100010011100100000000000000011001110001000000000111100010100000000001011100101000110001010101111100111111100101000000000000000000111110111001110011000000000000000000111011001010000010000000000000000000000101000100000000000000000011011110100000000100000000000000000000100001000000000000000000100000000010101101000000000000000000011100000000000000100000000000000000100000000001011001000000000001011100000000000100000000111011011011000110000000000100000000000000000010110010011011001100000000110110100000000000000000011111111111000000000000011011010001110101001101100000000001011110001010101100000000001100011000000000111010111000010110111110011000000000110110011001111000111111110000000000000010010000000000000000100000000000001111011001110001000110000000000000111000110100000000000000000101110010001110111000000000010110101000000000100000000010011111111010101000000000010000111101110101111111010101001110100000000100000000000000000010000110101000101111111000010110000100010000001000100000000000100000000000000000111110101101001000101001110000010111100000000010101111000000000111110111000001001100000000000000000000000000100000000000000000000001110001101100000000000; 
         #10 
        bram_addr_a2 = 6;
        weight_write = 1260'b110000000001100011000000000011000100100000000100000000000000000000000000100000000001001100000000100001001101100000000000000011110101111000000000001001011100000000001000001000000000000000000010011011001010010000000000011111100000110110100000000000000000000000000100000000010001000000000000000000000100000000001111000000000000111100010000000000100000000000000000000011011000000000000000000001111110010110010000000000010010110100000000000000000000000000000000000001011110000101111000000000000101000000000000110101111000000100000000000000000000011101001000000000010011110100000000100000000010001001000000000000100110001000111000000000111011000000000000111010011010111000100000000001010101100000000110101011000000000010001001000101011000000000000000000001111000001100101100000000111000111101101010000000000111111110000000000111001010000000000000000000000000000000011011001101100000000000010110001111010010000000000100011101000000000000000000111100101100000000000000000100000000100000000100000000010001111001101111100000000000000000101111100100000000000000001100000001001010111001010000000000000100000000000000000111101000000000000010011111100000000100000000100111010000000000001101111000010010100000000011000110011111111100000000000000000010101011100000000000000000;
         #10 
        bram_addr_a2 = 7;
        weight_write = 1260'b001000011100000000000111011000000000001001000100000000000000000110010011010001111110001100111110001100000000100000000111111010100000000000000000100000000100000000111001101010100111001010101100000000101001001000000000000000000100000000100000000000000000000000000001100100100010110000000000000000000010101000010110111000000000100000000011000100000000000000000000101111011010001110000000000100000000100000000000000000101101011101111001000000000000000000000000000000000000100000000000000000110101001000000000010111101000000100000000000011110001100000000000111001100000000000000000100000000100000000000000000101111110000110011000000000000100000000000000000101001100000000100000000000010011010100100000000000011100011100110101101111001100000000000000000101000001100000000111110001000000000001000000000000000000000110000000000100000000000000000001001001010110001101101100100000000000000000000000000100000000000000000100000000000000000000000000100000000010110111011111111010101001100000000001111110100000000110100110001011011000000000000000000001100110000000001100000000110110111100010001000000000000100100000000000000001011101001000100000000000010111010001000100000000000000000100000000111011111100000000000000000000000000100001010000000000110011011100111010010111111; 
         #10 
        bram_addr_a2 = 8;
        weight_write = 1260'b110000000100000000010000110100000000110100000000101011000000000100000000000110101101001011000000100001101001111100101000000011001110001000000000000100110111100000111111010001001100001010101010000001000001111000000000000000000001001001000111110000000000000000000000101010110100011000000000000000000100000000000000000000000000001111110100000000000000000000000000000100001000000000000000000011001011100000000111000111100000000111001101000000000010100100000000000000000000000111110000000000000010001000000000101110010000000001011000110000000000100000000000000000110001010000010001011011001010100110000000000000000011110001111000000000000011011000000000001011011010110100111100111011000011000000000000000000000000000111010111111000100001110000000000000001100111101111110101100101000000000111101000000000000000000001000000000001001111000000000000110000000000000111010011100000000000000000000000000010101011000000000001110001000000000000000000001011100000000000000000000000111101101110101100000000111011000100000000100000000000000000001100000100000000111111111010010101100000000111001111000000000000010010000000000000001000000000000110001000100000000000001011010011000000110010001011110000010111111011100000000000000000000011100110000000000000000000000011010100000000; 
         #10 
        bram_addr_a2 = 9;
        weight_write = 1260'b000111110000000000010101011100000000110100000010100110000000000010101001000100101101110011000000110100000000100000000000000110000000000000000000001110000100000000100000000010101100000000000100000000111010011000000000000000000000110010110010010000000000000000000100000000101111110000000000000000000001001100000000000000000000100000000001101101000000000000000000111011100100000000000000000100100011100000000011010111100000000100000000000000000100000000000000000100000000100000000000000000110110001000000000100000000000000110000000000000000000000000000000000000100000000000000000000100001101110010000000000000110000000111110000000000000011000000000000001010100100001010100000000000000000010101111110101011000000000100110101000101110100000000000000000100000000100010110110011001000000000000000111000000000000001001000000000010111010001110001100000000011010101000100110100000000100000000000000000100000000000000000000000000001110001100000000100000000100000000000000000010010000111101110001001011100000000000000000010110000000000000100000000000100010000000100100000001000110101100000000000000000000110110000000000000001110111100100000000000001111100000100100010100011101001000010100001000010100010000011000000000000000000000010011000000000100000000000000000011001000; 
        #10 
        bram_addr_a2 = 10;
        #10 
        bram_addr_a = 0;
        clause_write = 0;
	#10
bram_addr_a = 0;
clause_write = 182'b10100101110010000000000011011001110111110111101000000000000000000000000000000000000000011011110000000000000000000000000111001110010100111001110000000000000000;
#10
bram_addr_a = 1;
clause_write = 182'b11110100101111000000000111011111111100000000000000010000010000010000100000000000000000001111110000000000000000000011101111000110000100001000000000000000000000;
#10
bram_addr_a = 2;
clause_write = 182'b00010000100000001000000000010001100100000000000010100000000000000000000000000000000000000001000000000000000000000000000000000001000010011010010000000000000000;
#10
bram_addr_a = 3;
clause_write = 182'b11000101100001000001000010101000000000000000000000000000000000000000001000000000000000000000000000000000000000011000001100110110000010000100000000000000000000;
#10
bram_addr_a = 4;
clause_write = 182'b00010000000000000000000100011000000000000000000000000000000000001000100000000000100000000000000000000000100100000000000001000000000100001000010000000000000000;
#10
bram_addr_a = 5;
clause_write = 182'b11111111111110000000000111111000000000000000000000100000000000000000000000000000000000111111110000000111111111101111111100111101111111111111110000000000000000;
#10
bram_addr_a = 6;
clause_write = 182'b00000000100000000000000000000110110000000000001000010000000011000001100000000000000010010000000000000000000010100000000100001000000000000000000000000000000000;
#10
bram_addr_a = 7;
clause_write = 182'b11111111111111111111100111111100000000000000001111101111001100000000000000000000000000000000010000000000001111111111100000000000000011111111110000000000000000;
#10
bram_addr_a = 8;
clause_write = 182'b10000000000000000000000010011100000101100001100000000000100001000010000000000000100001100000000000000000000000000000000001001110010000010000010000000000000000;
#10
bram_addr_a = 9;
clause_write = 182'b00001000000000000000000000000000010010000000000000000000001000001000010000000000001101000000000000000000000000000000010000100000100011000010000000000000000000;
#10
bram_addr_a = 10;
clause_write = 182'b11111101111111000000000100000000000000000000000000000000000000000100001000000000000000011011100001111110100011111110111111101011111001000110000000000000000000;
#10
bram_addr_a = 11;
clause_write = 182'b11101111100000000000000100000000000000000000000000100001000010000100001000000000000001111110110001111111101101101111111100110001110011100010000000000000000000;
#10
bram_addr_a = 12;
clause_write = 182'b10000000000000000000000111111111110000000000000000000000000001110011111000111111111111111011110000000000001111111111111111111111111100000000000000000000000000;
#10
bram_addr_a = 13;
clause_write = 182'b11010000000000000000000111111000000000000000000000000011001000100010000000000111001111111111100000000000001111110011111000100000000000011001110000000000000000;
#10
bram_addr_a = 14;
clause_write = 182'b01000000011000000000000000000000000000000000000000100000000110001100011000000000000010000010010000000000000000101100001000100001000001100010000000000000000000;
#10
bram_addr_a = 15;
clause_write = 182'b11111111100000000000000110011011111111111100001000011000100001000010000000000000000111110111010000000000000000000000100111000100011100111001010000000000000000;
#10
bram_addr_a = 16;
clause_write = 182'b00000000000000000000000000000000000000000000000000000100001000000000000000000000000101001001000000000010000000101110010000000000000110000011110000000000000000;
#10
bram_addr_a = 17;
clause_write = 182'b11010101000000000000000010111100000000000000001000011001011100000000000000000000001110111111110000000000000011011111100100000000000000000000000000000000000000;
#10
bram_addr_a = 18;
clause_write = 182'b11100000000000000000000111111111111111111000000000000000000000000000000000111111111111111111110000000000000000011111111111111111111111111111110000000000000000;
#10
bram_addr_a = 19;
clause_write = 182'b11000111000000000000000111101000000000000000000000000001000110111011110000000000011110111111110000000000011111011111111100110001000000000000000000000000000000;
#10
bram_addr_a = 20;
clause_write = 182'b11111111111110000000000111111111111111111100001100011000110001000000000000000000000000111111110000000000000000000000100011000110001100011001110000000000000000;
#10
bram_addr_a = 21;
clause_write = 182'b01110011110111011100000101011000000000000000000001100000000000000000000000000000000000000001110000000010111110111001010000111001111011001001110000000000000000;
#10
bram_addr_a = 22;
clause_write = 182'b01000000000000000000000111111111100000000000000000000000000000000100001000111111111111111111110000000000001111111111111111111111111011110011000000000000000000;
#10
bram_addr_a = 23;
clause_write = 182'b00000000000101000000000000000001010000000000001000010000100000000000001000000000000000000000000000000000000010000000000000000000010000000000000000000000000000;
#10
bram_addr_a = 24;
clause_write = 182'b00000000000000000000000100010100101101000000001110000000000000000000000000000001011100001100100000000000000000000000000000000001101110110101110000000000000000;
#10
bram_addr_a = 25;
clause_write = 182'b00000000000000000000000000001000100000000000001000000000000000000000000000001011010001000100100000000000000000000110100001000010010111100101010000000000000000;
#10
bram_addr_a = 26;
clause_write = 182'b11111111111111110000000110000000000000000000000000000000000000000000001000000000000000000011010000111111111111111111111111111111111111110111000000000000000000;
#10
bram_addr_a = 27;
clause_write = 182'b00000100000000000000000000000000100000011000000010000000000000000000000000000000000100100000000000000000000000000000000000000000010111010010000000000000000000;
#10
bram_addr_a = 28;
clause_write = 182'b00000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
bram_addr_a = 29;
clause_write = 182'b00100011000010000010000001000010000000000000000000000000000000000110000000000000000000000000000000000000000000010100000000000000010000000000000000000000000000;
#10
bram_addr_a = 30;
clause_write = 182'b11000000000000000000000111011111101100000000000000000000001000110011100001111111111111111111100000000000000000011011111111100100000000000000000000000000000000;
#10
bram_addr_a = 31;
clause_write = 182'b00000100000000000000000000000000000000010000000000000000000000001000000000000000010000000000000000000000000000000000011100010000100000000000000000000000000000;
#10
bram_addr_a = 32;
clause_write = 182'b10000000000000000000000111111111000000000000000000000000000000000000001011111111111111111111110000000000111111111111111111111111111111110111000000000000000000;
#10
bram_addr_a = 33;
clause_write = 182'b00011000000000000000000101000010000110000000000000000000000000000011011000000001000000000000000000000000000000000000000000100101100000000000000000000000000000;
#10
bram_addr_a = 34;
clause_write = 182'b10011110111101000000000001011111000000000000000000100001000010001100001000000000000000000001000000000000011010111001111100111000010011100111000000000000000000;
#10
bram_addr_a = 35;
clause_write = 182'b11111111111111110000000111110111111111000000001100011000110001000000000000000000000000000111110000000000000000011111100011000110011100111011110000000000000000;
#10
bram_addr_a = 36;
clause_write = 182'b11111111110100000000000111011101110111111000000000000000000000000001000000000000000000001110100000000000000000000001101111011111100100000000000000000000000000;
#10
bram_addr_a = 37;
clause_write = 182'b00000000000000000000000111111111111101000000000000000000000000000010000111111111111111111111110000000000000000011111111111111111111111111000110000000000000000;
#10
bram_addr_a = 38;
clause_write = 182'b11010110011111000000000110000000000000000000000000100100010000100001000000000000000000000111000000000010011000000110000000000000000000010000000000000000000000;
#10
bram_addr_a = 39;
clause_write = 182'b10111111101110100000000101000111110000000000000011001100010001011001111000000000000000000011010000000000000111100011000000000000000000000000000000000000000000;
#10
bram_addr_a = 40;
clause_write = 182'b11111111111110000000000000000000000000000000000000000001000000000000000000000000000000011111110011111111011111111111111110111101111011110111100000000000000000;
#10
bram_addr_a = 41;
clause_write = 182'b00000000000000000000000000000000000011000000000000000000000000000100000000001000000000000000000000000000000000000000010000010000110001000110000000000000000000;
#10
bram_addr_a = 42;
clause_write = 182'b10111111001000000000000010100000111100000000000000000011000100011000100000000000000011100110000000000000000000001101101000010000100010000100000000000000000000;
#10
bram_addr_a = 43;
clause_write = 182'b11000000000000000000000000000101011100000000000000000000000000000100110000010000000010100111100000000000000000101010000110101101011011000100000000000000000000;
#10
bram_addr_a = 44;
clause_write = 182'b10000000000000000000000101111111000000000000000000000000000000111011111001111111111111101111110000000000001011111110111111111111111100000000000000000000000000;
#10
bram_addr_a = 45;
clause_write = 182'b11111111100000000000000111111100000000000000000100011000110001111101111000000000001111111111010000000000111111111111100000000010000000000000000000000000000000;
#10
bram_addr_a = 46;
clause_write = 182'b00000010100111000000000110000000000000000000000000000000000000000000100000000000000000001111100000000000101101011010111010011010000100001000000000000000000000;
#10
bram_addr_a = 47;
clause_write = 182'b00000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000100000000101000000000110010000001000000100000000000000000000000000;
#10
bram_addr_a = 48;
clause_write = 182'b00000100000010000000000000000000110000000000000000000000000000000000000000000000000000100000000000000000000101000000011000000100000110000101010000000000000000;
#10
bram_addr_a = 49;
clause_write = 182'b00110110000000000000000001000000000000000000000000000000000001011111111000000000000000111110110000000110101101111011110000100000000000000000000000000000000000;
#10
bram_addr_a = 50;
clause_write = 182'b01011110111101000000000111000000000000000000000001000100001000010000100000000000000000000111110000000001100110011100100000000000000100001100000000000000000000;
#10
bram_addr_a = 51;
clause_write = 182'b00000101000110010110000000010100111010000000000000000000100000000000000000000000000000000000000000000000000000000000011101000000001000100000010000000000000000;
#10
bram_addr_a = 52;
clause_write = 182'b11000000000000000000000111110000000000000000000000000000000000000000001000111111111111111111110000001111111111111111111111111111111111111111100000000000000000;
#10
bram_addr_a = 53;
clause_write = 182'b11110111111000000000000111010100111100000000000000000000000000000000000000000000000001111011110000000000000001110100101111001110101101111011110000000000000000;
#10
bram_addr_a = 54;
clause_write = 182'b11111111111111100000000111111111111111111000001100000000000000000000000000000000000000001111010000000000000000000000100011001111111111111111110000000000000000;
#10
bram_addr_a = 55;
clause_write = 182'b00000000000000000000000000000000000000000000000000100000000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
bram_addr_a = 56;
clause_write = 182'b00000000010000000000000000000000100100000000000110000100001000100000000000000000000001001100000000000000000011010000000001000010001000000000110000000000000000;
#10
bram_addr_a = 57;
clause_write = 182'b11100000000000000000000111110000000000000000000000000000000010000100001000000111111110100111110000001111111111111111111110111101011011100111000000000000000000;
#10
bram_addr_a = 58;
clause_write = 182'b11111000000000000000000110011011111101111111000000000000000000000010000000000011101101011101110000000000000000000000101111010111101101011001110000000000000000;
#10
bram_addr_a = 59;
clause_write = 182'b11111111100011000000000111111100000000000000000001101011000100110001100000000000000000001111010000000001100111100110100000000000000000000000000000000000000000;
#10
bram_addr_a = 60;
clause_write = 182'b11100000000000000000000111111110111000000000000000000000000110111111000000010111101110111111100000000000000000111110111111110111100000000000000000000000000000;
#10
bram_addr_a = 61;
clause_write = 182'b00111110000000000000000011011011111100000000001011111100000010000100010000000000100001111111010000000000000000010111100000000000000000000100000000000000000000;
#10
bram_addr_a = 62;
clause_write = 182'b11111011000000000000000111101101101111110000000010001000100000000000000000000000001011111111110000000000000000000111000000000010000001111111110000000000000000;
#10
bram_addr_a = 63;
clause_write = 182'b01011111111111011111010111111111001100000000001111011000000000000000000000000000000000000000000000000000000001111110100000000010101011111110110000000000000000;
#10
bram_addr_a = 64;
clause_write = 182'b00001000000000000000000001000000000000000000000000000000000000000001000000000010000000000000000000000000100010000000000001000010000100001000010000000000000000;
#10
bram_addr_a = 65;
clause_write = 182'b11100000000000000000000111101111111111111110000000000000100000000000000000011111111111111111110000000000000000000001111010001110010100110001110000000000000000;
#10
bram_addr_a = 66;
clause_write = 182'b11111111111111111111100111111111111111000000001000010000100000000000000000000000000000000000010000000000000000011111100111001110011101111111110000000000000000;
#10
bram_addr_a = 67;
clause_write = 182'b11111000000000000000000000000000000000000000000000000001000000000000000000000000011111110011100010110111110111101111110000101001000001000101100000000000000000;
#10
bram_addr_a = 68;
clause_write = 182'b11111111111101101100000111111110000000000000000000000000000000000000000000000000000000000111110000000001111110110111111111111111111111010111110000000000000000;
#10
bram_addr_a = 69;
clause_write = 182'b00000000000110000000100000000000000100000000000010000000000000010000000000000000000000000000000000000000000000000001000000000000000010000100000000000000000000;
#10
bram_addr_a = 70;
clause_write = 182'b11101111010000000000000001111111011111011110001000000000000000000000000000000000001111100111110000000000000000000001100110011011111111111111110000000000000000;
#10
bram_addr_a = 71;
clause_write = 182'b10011111111010001110000111101111000000000000001100000011000000000000000000000000000000000001110000000000000001101111100000000000000010111110110000000000000000;
#10
bram_addr_a = 72;
clause_write = 182'b00010100000000000111000100010000000000000000000000000000000100000000000000000000000000000000000000000000000000111000001011100001000010000100000000000000000000;
#10
bram_addr_a = 73;
clause_write = 182'b00000100000000000000000000000000000000000000000100010000000001000000001000000000000001100000000000000100000000000001000000000110000000000000000000000000000000;
#10
bram_addr_a = 74;
clause_write = 182'b00000011000000000000000000011000000000000000000010000100000010000000000000000000000000001000000000000000100000000000100001010000000000100100000000000000000000;
#10
bram_addr_a = 75;
clause_write = 182'b00000000000000000000000000000000000000000010001011000000000000000000000000000000000000000000000000000000000000000000000000000001100010001111100000000000000000;
#10
bram_addr_a = 76;
clause_write = 182'b01011110000000000000000111111111110111111101100000000000000000000011000000000000000000110111110000000000000000000000000001000000000100000000110000000000000000;
#10
bram_addr_a = 77;
clause_write = 182'b00000000000000000000000000000000000000000000000010000000000010000010100000000000100000000000000000000000000000000000000000000000010000000000000000000000000000;
#10
bram_addr_a = 78;
clause_write = 182'b11111111111101111111000111111000000000000000001000011001011100000000000000000000000000000000010000000011111111111101100000000000000000000111110000000000000000;
#10
bram_addr_a = 79;
clause_write = 182'b00000000000000000000000100001000000000000000000000100000000000000000000000000011100000000000000000000000010110000010110000000001000010001111000000000000000000;
#10
bram_addr_a = 80;
clause_write = 182'b00000000000000000000000100111010001111111101010000000000000000000000000011101111111111101011110000000000000000000000011111110111110101111111110000000000000000;
#10
bram_addr_a = 81;
clause_write = 182'b00000000000000000000000000000000000000000000000000100000000000000000000000000110000011100000010000000000000111100100110000000001000001111101000000000000000000;
#10
bram_addr_a = 82;
clause_write = 182'b11111000000000000000000111110000000000000000000000000000000000000000001000001111111111111111110000000111111111111111111111111111111111111111100000000000000000;
#10
bram_addr_a = 83;
clause_write = 182'b11111000000000000000000111111111111111111000000000000000000000000000000000001111111111111111110000000000000000001111111111111111111111111111110000000000000000;
#10
bram_addr_a = 84;
clause_write = 182'b11100000000000000000000111111111101111111110000000000000000000000011000000011111111011111111110000000000000000000000001111111111111100111000110000000000000000;
#10
bram_addr_a = 85;
clause_write = 182'b10001000000010000000000000000000100101000000000000000000000000000011110000000000000000000000000000000000000000000000000010101001000000000000000000000000000000;
#10
bram_addr_a = 86;
clause_write = 182'b11101000000000000000000111111111100000000000000111001111111100111011110000000001111111111111110000000000000000011111100000000000000000000000000000000000000000;
#10
bram_addr_a = 87;
clause_write = 182'b00100000000000000000000111001000000000000000000000000000001000000001110000110100100100001001000000000000000111110100100110000010000000000000000000000000000000;
#10
bram_addr_a = 88;
clause_write = 182'b00000000000000000000000000000000000000000000000000000000010000000010000000000100000000000000000000000000001000000000000010000100000000010000110000000000000000;
#10
bram_addr_a = 89;
clause_write = 182'b00000010000000000000000000000010000000000000000001000010000010000100001000000000000000000010000000000000110000000000010000010000010000000101000000000000000000;
#10
bram_addr_a = 90;
clause_write = 182'b11111111111111111111100111110000000000000000000000100000000000000000000000000000000000000000010000001111111111111111111110111101111111111111110000000000000000;
#10
bram_addr_a = 91;
clause_write = 182'b11111101101000000000000111111011111100000000000001110111101110101101110000000000000000011001100000000000000001111111000000000000000000000000000000000000000000;
#10
bram_addr_a = 92;
clause_write = 182'b11000000000000000000000111001111110110000000000000000000000001110001110000111110110111111110110000000000000000001111101011011111111100001000000000000000000000;
#10
bram_addr_a = 93;
clause_write = 182'b11111100000000000000000111111011111111110000000000000000100001000010000000000000101110111101110000000000000000001111111111011110011100111001100000000000000000;
#10
bram_addr_a = 94;
clause_write = 182'b00000000000000000000000110110100000000000000000000000000000000000000001110111101110111111101110000000000011010110110111110001100111011111110000000000000000000;
#10
bram_addr_a = 95;
clause_write = 182'b11111111111010000000000111100111101111100000000100011000110001000000000000000000000000111110110000000000000000011110100001000010011100111011100000000000000000;
#10
bram_addr_a = 96;
clause_write = 182'b10110101101010110000000000100101011011100000000000000000000000000010000000000000000000000011110000000000000000000100001111111100000100000000000000000000000000;
#10
bram_addr_a = 97;
clause_write = 182'b01000000000000000000000111111011101100000000000000000000000000000011110000111111111111111111100000000000000000000001111111110111111111111000000000000000000000;
#10
bram_addr_a = 98;
clause_write = 182'b00101011010000000000000000000010100000000000000000000001001000000000000000000000000100000100000000000000000000000000000000000000000010000001100000000000000000;
#10
bram_addr_a = 99;
clause_write = 182'b11111010110110000000000111000011000000000000000100001111000010000000000000000000000000111101110000000000000111011101100000000000000011110000100000000000000000;
#10
bram_addr_a = 100;
clause_write = 182'b00111111111111110000000010001110001000000000000001100100110100010010000000000000000000000000010000000000000001000110010000000000000000001001110000000000000000;
#10
bram_addr_a = 101;
clause_write = 182'b11111111110000000000000110101111111111110000000000000000000001110000000000000000000011111111110000000000000000000001111111001110000100001000000000000000000000;
#10
bram_addr_a = 102;
clause_write = 182'b11111111111111111110000111000000000000000000000001100001000000000000000000000000000000000000110000011111111111111111111100111001111011111111110000000000000000;
#10
bram_addr_a = 103;
clause_write = 182'b11111111111111111111000111100000000000000000000111100011000000000000000000000000000000000000000000001111111111111111100000000001111010111111110000000000000000;
#10
bram_addr_a = 104;
clause_write = 182'b00000010100000010011100001000000000000000000000000100010000000010000100000000000000000000000000000000000000110000001000000100000000000000100000000000000000000;
#10
bram_addr_a = 105;
clause_write = 182'b01010000000000000000000111000011110100100000000000011000010001000010000000000001101101011100100000000000000000010000100011001010011100001001000000000000000000;
#10
bram_addr_a = 106;
clause_write = 182'b01001100010000000000000000000000000000000000001000000000100000100000111000000000000010110000000000000101000100011010100000000010001000000000000000000000000000;
#10
bram_addr_a = 107;
clause_write = 182'b01000000100000000000000000100000000000000000000000000000000000000001100000000000000010001010010000000001100000100000010000010001111110000000000000000000000000;
#10
bram_addr_a = 108;
clause_write = 182'b11101111111110000000000111111100000000000000000000000000000000000000001000000000000000111111110000000001111111111111111111111111111011110111000000000000000000;
#10
bram_addr_a = 109;
clause_write = 182'b00110000000000000000000000111010111011000000000011000100010001000010000000000011111111111111010000000000000000000001100000000000000100011001010000000000000000;
#10
bram_addr_a = 110;
clause_write = 182'b11001011011110111110000111111101000000000000001000111101111101110000000000000000000000000000010000000000000001111101100000000000000000000011110000000000000000;
#10
bram_addr_a = 111;
clause_write = 182'b11111000000000000000000111111111111111100000000000000000100001100011000000000111111111111111110000000000000000001111111111011110011100011000010000000000000000;
#10
bram_addr_a = 112;
clause_write = 182'b00000000000000001000000000000000000001100000000001000000000000000000000000000000000000000000000000000000000000000000010000010001100000100000100000000000000000;
#10
bram_addr_a = 113;
clause_write = 182'b00111100111000100000000000001111100000000000000010001000111000000001000000000000000000000000000000000000001100010110000000000010001100001000110000000000000000;
#10
bram_addr_a = 114;
clause_write = 182'b00000010000000000000000000000000010010000000000011000000000000000000000000000000010000000000000000000000000000000000000000000001110010010000110000000000000000;
#10
bram_addr_a = 115;
clause_write = 182'b00101011010000000000000100000000000000000000000000000000000000000100011000000000001011000010110000011110000101111101110111010110111001100000000000000000000000;
#10
bram_addr_a = 116;
clause_write = 182'b11100000000000000000000011111110111111000000001100000000000000000000000000000101111111111110100000000000000000000000000001000110011111111111100000000000000000;
#10
bram_addr_a = 117;
clause_write = 182'b00000000000000000000000010000000000000000000000000001000010001000010000000000110100001000000010000000000000011000010000011000010001100011000100000000000000000;
#10
bram_addr_a = 118;
clause_write = 182'b00000000000000000000000111111000000000000000000000000000000000000000001111111110101111111111000000000000111111111111111111111111111011110111000000000000000000;
#10
bram_addr_a = 119;
clause_write = 182'b00000000000000000000000100000000000000000000000000000000000000000010000000000010000000000010000000000011000000000000010001000100000100010000000000000000000000;
#10
bram_addr_a = 120;
clause_write = 182'b00010100000111000000000000000000000000000000000000100010001000000000110000000000000000000011110000010101101111011000001000000000000010000000000000000000000000;
#10
bram_addr_a = 121;
clause_write = 182'b10100000000000000000000000111000000000000000000110000000000000000000001000000000000011110011100000000001101001111001000000000001110000000100000000000000000000;
#10
bram_addr_a = 122;
clause_write = 182'b00000000110100000000000000000000000100000000001110100001000100010001000000000000000000011000000000000000000001100000000000000000000000001000110000000000000000;
#10
bram_addr_a = 123;
clause_write = 182'b00101100011100001111000011111100101110000000000000000010001000000000000000000000000000000000000000000000000000000111011000000000000000000001100000000000000000;
#10
bram_addr_a = 124;
clause_write = 182'b11101100000110000000000111111110111111111100001000000000000000000000000000000000000001101110110000000000000000000001100110111111110111110110110000000000000000;
#10
bram_addr_a = 125;
clause_write = 182'b00110011110000000000000111100100010010000000001110010100001000110001000000000000000001110010110000000000000000101100100000000010000100010000100000000000000000;
#10
bram_addr_a = 126;
clause_write = 182'b11111111111111111100000111000000000000000000001011111101011000000000000000000000000000000001110000000000011101111111100000000000000000001111110000000000000000;
#10
bram_addr_a = 127;
clause_write = 182'b11100011000000000000000110111100000000000000000000000001000110000000100000000000001011100001100000000011000011010000010010111000010010000100000000000000000000;
#10
bram_addr_a = 128;
clause_write = 182'b11111110000000000000000100000000000000000000000001100000000000000000000000000000011011111111110000011111111111001111110000100001100011100111110000000000000000;
#10
bram_addr_a = 129;
clause_write = 182'b11110000000000000000000111111111100000000000000000000111011110111111001000000111111111111011110000000000001111011111110000000000000000000000000000000000000000;
#10
bram_addr_a = 130;
clause_write = 182'b11000000000000000000000110101100000000000000000000000000000000000100011000111111111111111111110000000001110111110111010101111111000110100110000000000000000000;
#10
bram_addr_a = 131;
clause_write = 182'b10000000000000000000000111111111000000000000000000000000000001111111011001111101111111111111010000000000000011111111111111111111000000000000000000000000000000;
#10
bram_addr_a = 132;
clause_write = 182'b11111111111111111111100111111111100000000000000000000000000000000000000000000000000000000000110000000000011111111111111111111111111111111111110000000000000000;
#10
bram_addr_a = 133;
clause_write = 182'b00000001000100000000000000000010000000100000000100000100000000001000000000000000000000000110000000000000000000000000000001000000100000000000000000000000000000;
#10
bram_addr_a = 134;
clause_write = 182'b10001010000000000000000011000000000000000000000000010000010000110000101000000000010001001011100000000000111011101011000000000000000100000000000000000000000000;
#10
bram_addr_a = 135;
clause_write = 182'b01111110000000000000000000100100000000000000000000001111011110000000000000000000111110110011100000000000000000000011100000000000000000000101110000000000000000;
#10
bram_addr_a = 136;
clause_write = 182'b11100000000000000000000111111111100000000000000000000000011001111111111000011111111111111111110000000000000011111101110111111010000000000000000000000000000000;
#10
bram_addr_a = 137;
clause_write = 182'b00101000011010000000000100001100000000000000000001100001011000000110001000000000000000001110010000000000100110001001000000000000000000000000000000000000000000;
#10
bram_addr_a = 138;
clause_write = 182'b00000000000000000010000000000000000000000000000100000000000001000000000000000000000000000000000000000000010000000000100001000000000100001000100000000000000000;
#10
bram_addr_a = 139;
clause_write = 182'b00000000100000000000000000000000001000000000000000000000101000010000010000000000000010000000000000000000000000100000001000001010000100000000000000000000000000;

                #10
        bram_addr_a = 140;
        end
//        always @(posedge output_params[4]) begin
//        count = count + 1;
//        #10
//        prst[1] = 1'b1;
//        #10 prst[1] = 1'b0;
//        #10
//             if(count == 1)begin
////         //number 1
//         total_img = 512'b00000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000;     
//        end
//        else if(count == 2)begin
//         //number 2
//         total_img = 512'b10000000000000000000011111000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001111010000000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000011110000000000000111111111111111000000000000111111111111111100000000000001000000111111;     
//        end
//        else if(count == 3)begin
//         //number 3
//         total_img = 512'b00000000000000000110000000000000000000000000011100000000000000000000000000111100000000000000000000000001111100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000000100000000000000000000000000110000000110000000000000000011000000111000000000000000001100001111000000000000000000111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000000011100011100000000000000000011000000110000000000000000001100000110000000000000000000110000010000;     
//        end
//        else if(count == 4)begin
//         //number 4
//         total_img = 512'b11000000000000000111111111111100000000000000011100000111100000000000000000110000111100000000000000000011100011100000000000000000001110011110000000000000000000110011110000000000000000000011001110000000000000000000001101110000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000000111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111111111111000000000000000011111111111;     
//        end
//        else if(count == 5)begin
//         //number 5
//         total_img = 512'b10000000000000001100000000011000000000000000110000000001000000000000000011100000000000000000000000000111100000000000000000000000001111111110000000000000000000001111111000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000010001111100000000000000001111111111100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//         total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111110000000000000000011110000111100000000000000001110000000110000000000000001110000000011000000000000000110000000001;     
//        end
//        else if(count == 6)begin
//         //number 6
//         total_img = 512'b00000000000000111110111111110000000000000011101111111111000000000000001111111110111100000000000000111111100011110000000000000011111100001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000001111110000000000000000000100111110000000000000000000111111110000000000000000000111111110000000000000000000011111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111110000000000000000011111111111100000000000000011111111111110000000000000001111101111111;     
//        end
//        else if(count == 7)begin
//         //number 7
//         total_img = 512'b00000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000001111000000000000011111111111111111100000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000;     
//        end
//        else if(count == 8)begin
//         //number 8
//         total_img = 512'b00000000000000000000111111100000000000000000000011111100000000000000000000001111100000000000000000000001111110000000000000000000001111111000000000000000000001111111100000000000000000001111001110000000000000000001111000011100000000000000000111000111110000000000000000111111111110000000000000000011111111110000000000000000001110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111110000000000000000000001111111000000000000000000001111011100000000000000000001111001110000000000000000000111000110000000000000000000011101111;     
//        end
//        else if(count == 9)begin
//         //number 9
//         total_img = 512'b00000000000000000011100000000000000000000000001110011111000000000000000000110011111100000000000000000111011111111000000000000000011111100011100000000000000001111000001100000000000000001111000001110000000000000000111000011110000000000000000111100111110000000000000000011111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000;     
//        end
always @(posedge opm) begin
    label = (img_count)/996;
    if(label == calc_label)success = success + 1;
    else fail = fail + 1;
    #10 prst[1] = 1'b1;
    #10 prst[1] = 1'b0;
    #10 load_next_chunk();
    #10 load_next_chunk();
end
always @(posedge clk) begin
calc_label = output_params[3:0];
opm <= output_params[4];
end
reg [511:0] total_img;
integer fd, r;
reg [1024*8:1] line; // buffer for each line
reg [783:0] bits784;
integer j;
integer cycle_count = 0;

initial begin
    fd = $fopen("10ktest.hex","r");
    if (fd == 0) begin
        $display("Error: could not open file");
        $finish;
    end
end

task load_next_chunk;
        begin
            if (cycle_count == 0) begin
                // read one image = 784 ASCII chars
                for (j=0; j<784; j=j+1) begin
                    r = $fgetc(fd);
                    if (r == "0")
                        bits784[783-j] = 1'b0;
                    else if (r == "1")
                        bits784[783-j] = 1'b1;
                    else
                        j = j - 1; // skip newline or junk
                end
                // chunk 1 = lower 512
                total_img = bits784[511:0];
                cycle_count = 1;
            end
            else begin
                // chunk 2 = upper 271 + padding
                total_img = {241'b0, bits784[783:512]};
                cycle_count = 0;
                img_count = img_count + 1;
            end
        end
    endtask
        
endmodule
